module can_defines