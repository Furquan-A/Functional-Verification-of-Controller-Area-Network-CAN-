class can_bus_model extends 