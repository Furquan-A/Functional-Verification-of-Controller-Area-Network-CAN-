class env extends uvm_env;