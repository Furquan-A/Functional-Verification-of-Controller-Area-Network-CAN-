class can_frame_sequence extends uvm_items ;
