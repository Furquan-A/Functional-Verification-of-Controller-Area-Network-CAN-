class can_stress_test extends uvm_tests;
