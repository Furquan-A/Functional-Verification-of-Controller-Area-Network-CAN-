class can_basic_test extends uvm_tests;
