class can_base_test extends uvm_test;