class can_driver extends uvm_componen