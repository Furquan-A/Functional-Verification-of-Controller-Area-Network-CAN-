class can_transactions extends uvm_transactions;