class can_virtual_sequences extends uvm_items;