class can_bit_timing_sva extends 