class can_frame_format_sva extends 