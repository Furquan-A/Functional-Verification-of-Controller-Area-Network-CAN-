class can_coverage extends uvm_items ;