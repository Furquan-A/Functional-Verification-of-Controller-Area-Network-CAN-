class reg_monitor extends uvm_component;