class can_config extends uvm_items;