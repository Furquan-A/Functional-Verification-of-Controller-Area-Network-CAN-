class can_sequence extends uvm_sequencer ;