class reg_seq extends uvm_items;