class can_scoreboard extends uvm_scoreboard;