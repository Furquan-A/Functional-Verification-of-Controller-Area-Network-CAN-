class reg_driver extends uvm_component;