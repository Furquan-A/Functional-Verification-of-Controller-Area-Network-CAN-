class can_stuff_rule_sva extends