class can_monitor extends uvm_component;