class can_base_seq extends uvm_items;