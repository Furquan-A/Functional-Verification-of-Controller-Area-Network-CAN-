class reg_sequencer extends uvm_components;