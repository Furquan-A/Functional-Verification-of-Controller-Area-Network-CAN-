class reg_agent extends uvm_component;