class can_virtual_sequencer extends 