class can_error_test extends uvm_tests;

